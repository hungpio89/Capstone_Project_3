library verilog;
use verilog.vl_types.all;
entity Thesis_Project_vlg_vec_tst is
end Thesis_Project_vlg_vec_tst;
