library verilog;
use verilog.vl_types.all;
entity or_1bit_vlg_vec_tst is
end or_1bit_vlg_vec_tst;
