module apb_interface										// & register block 
(
	// INPUT LOGIC CONFIGURATION
	//------------------CPU INPUT------------------------//
	input logic						PCLK,
	input logic						PRESETn,
	//---------------------------------------------------//
	
	//-----------------APB INTERFACE---------------------//
	input logic						transfer,			// correct address index or not (PSEL & PADDR[11:8])
	input logic 					PENABLE,
	input logic						PWRITE,
	
	input reg	 [   7 :   0] 	PADDR,
	input reg  	 [   7 :   0] 	PWDATA,				// reference is 16 bit, currently use 8 bit (know reason why use 16 -> CONFIGURATION OF UART 8 bits or 16 bits send each)
	
	
//	reg [  7 :  0] state;						//		0x004				  4			 RW				0x0				[3] RX buffer overrun, write 1 to clear.
//														//																					[2] TX buffer overrun, write 1 to clear.
//														//																					[1] RX buffer full, read-only.
//														//																					[0] TX buffer full, read-only
//														
//	reg [  7 :  0] ctrl;							//		0x008 			  7			 RW 				0x00 				[6] High-speed test mode for TX only.
//														//																					[5] RX overrun interrupt enable.
//														//																					[4] TX overrun interrupt enable.
//														//																					[3] RX interrupt enable.
//														//																					[2] TX interrupt enable.
//														//																					[1] RX enable.
//														//																					[0] TX enable
//					
	input reg	 [   3 :   0]  state_i,
	input reg	 [   6 :   0]  ctrl_i,
	//---------------------------------------------------//
	
	//------------------UART RETURN----------------------//
	input reg	 [	  7 :   0]	read_data,
	//---------------------------------------------------//
	
	//-------------------USER INPUT----------------------//
	input logic  [  19 :   0] 	desired_baud_rate,
	
	input logic 					TXdone, 
	input logic 					RXdone,
	
	input logic 					error_tx_detect, 
	input logic 					error_rx_detect,
	//---------------------------------------------------//
	
	//OUTPUT LOGIC ASSIGNMENT
	//--------------APB INTERFACE RETURN-----------------//
	output logic 					rx_buffer_overrun, 
	output logic 					tx_buffer_overrun,
	output logic 					uart_run_flag,		// to control the TX and RX operation (only active in case transmit or receive data)
	output logic					PREADY,				// used by Transmitter & Receiver block
	output logic [  12 :   0]	cd,
	output logic 					clk_div16,
	output reg 	 [	  3 :   0]  state,				
	output reg 	 [	  6 :   0]	ctrl,
	output reg 	 [   7 :   0] 	write_data,			// reference is 16 bit, currently use 8 bits
	
	output reg	 [  31 :   0] 	PRDATA
	//---------------------------------------------------//
);
	// Local signal define
	
	// Logic
	logic 							div16;
	logic			[  12 :   0]	actual_cd;	
	logic 		[   7 :   0] 	uart_data_mid;
	
	// Register
	reg			[   6 :   0] 	ctrl_mid;
	reg			[   7 :   0] 	base_offset; 	
	
	// Local signal assignment for PADDR
	genvar i;
	generate 
		for (i = 0; i < 8; i = i + 1) begin: offset_assignment
			assign base_offset[i] = PADDR[i];
		end
	endgenerate
	
	// Local signal assignment for ctrl
	genvar j;
	generate 
		for (j = 0; j < 2; j = j + 1) begin: ctrl_assignment
			assign ctrl_mid[j] = ctrl_i[j];
		end
			assign ctrl_mid[2] = error_tx_detect;
			assign ctrl_mid[3] = error_rx_detect;
		for (j = 4; j < 7; j = j + 1) begin: conn_ctrl_assignment
			assign ctrl_mid[j] = ctrl_i[j];
		end
	endgenerate
	
baud_rate_divisor 				BAUD_RATE_DIVISOR_BLOCK
(
	// INPUT LOGIC CONFIGURATION
										.clk					(PCLK),
										.rst_n				(PRESETn),
	 
	// OUTPUT LOGIC CONFIGURATION
										.clk_out				(clk_div16)
);
	
	// always loop for define cd for clock divisor counter
	always @(desired_baud_rate) begin	
		actual_cd = 13'd0;
		case(desired_baud_rate)
			20'd600   : actual_cd = 13'd5208;
			20'd4800	 : actual_cd = 13'd651;
			20'd9600	 : actual_cd = 13'd325;
			20'd19200 : actual_cd = 13'd162;
			20'd28800 : actual_cd = 13'd108;
			20'd38400 : actual_cd = 13'd81;
			20'd57600 : actual_cd = 13'd54;
			20'd115200: actual_cd = 13'd27;
			20'd230400: actual_cd = 13'd13;
			20'd460800: actual_cd = 13'd6;
			20'd921600: actual_cd = 13'd3;					// Maximum baudrate for normal UART
			default   :	actual_cd = 13'd325;				// default 9600
		endcase
	end
	
	// APB Interface
	always @(posedge PCLK or negedge PRESETn) begin
		if (!PRESETn) begin										// RESETn operation (reset all registers)
			uart_data_mid 	<= 8'b0;
			state 			<= 4'b0;
			ctrl				<= 7'b0;								// 7 bits if related to Docs
			PREADY			<= 1'b0;
			uart_run_flag  <= 1'b0;
		end 
		else begin
			uart_run_flag  <= 1'b0;
			PREADY			<= 1'b0;
			if (transfer && PENABLE) begin
				if (PWRITE) begin										// WRITING MODE
					case (base_offset)
					// Base Offset
						8'h0: begin
							ctrl		<= ctrl_mid;								// write 1 to ctrl[0]	// custom write only
							PREADY	<= 1'b1;
						end
						8'h4: begin
							rx_buffer_overrun <= state_i[3];
							tx_buffer_overrun <= state_i[2];
							state[3:0]			<= state_i[3:0];
							PREADY				<= 1'b1;
						end
						8'h8: begin 											// this process is for set up clock (custom from PCLK)
							for (int l = 0; l < 13; l = l + 1) begin: cd_assignment
								cd[l]	<= actual_cd[l];
							end
							PREADY	<= 1'b1;
						end
						default: begin
							uart_run_flag  <= 1'b1;
							uart_data_mid 	<= PWDATA[  7 :  0];
							if (TXdone) begin
								PREADY	<= 1'b1;
							end
						end
					endcase
				end 
				else if (!PWRITE) begin												// READING MODE
					case (base_offset)
						8'h0: begin 
							PRDATA 		<= {28'b0, state};
							PREADY		<= 1'b1;
						end
						8'h4: begin 
							ctrl 			<= ctrl_mid;
							PRDATA		<= {25'b0, ctrl_mid};
							PREADY		<= 1'b1;
						end	
						8'h8: begin
							PRDATA		<= {19'b0, actual_cd};
							PREADY		<= 1'b1;
						end
						default: begin
							uart_run_flag <= 1'b1;
							PRDATA 		  <= {24'b0, read_data};
							if (RXdone) begin
								PREADY	<= 1'b1;
							end
						end
					endcase
				end
			end
			else
				PREADY	<= 1'b0;
		end
	end
	
	// Local signal assignment for write_data
	genvar k;
	generate 
		for (k = 0; k < 8; k = k + 1) begin: data_write_assignment
			assign write_data[k] = uart_data_mid[k];
		end
	endgenerate
	
	
endmodule
