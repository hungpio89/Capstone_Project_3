library verilog;
use verilog.vl_types.all;
entity AHB_SLAVE_vlg_vec_tst is
end AHB_SLAVE_vlg_vec_tst;
