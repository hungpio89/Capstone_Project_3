library verilog;
use verilog.vl_types.all;
entity fifo_read_memory_vlg_vec_tst is
end fifo_read_memory_vlg_vec_tst;
