module Thesis_Project ();


endmodule
