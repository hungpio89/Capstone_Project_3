library verilog;
use verilog.vl_types.all;
entity pipeline_riscv_mod2_vlg_vec_tst is
end pipeline_riscv_mod2_vlg_vec_tst;
