library verilog;
use verilog.vl_types.all;
entity test_ver5 is
    port(
        PCLK            : in     vl_logic;
        UARTCLK         : in     vl_logic;
        PRESETn         : in     vl_logic;
        desired_baud_rate: in     vl_logic_vector(19 downto 0);
        UART_RXD        : in     vl_logic;
        parity_bit_mode : in     vl_logic;
        stop_bit_twice  : in     vl_logic;
        uart_mode_clk_sel: in     vl_logic;
        number_data_receive: in     vl_logic_vector(3 downto 0);
        ctrl_i          : in     vl_logic_vector(6 downto 0);
        state_isr       : in     vl_logic_vector(1 downto 0);
        PSEL            : in     vl_logic;
        PENABLE         : in     vl_logic;
        PWRITE          : in     vl_logic;
        PADDR           : in     vl_logic_vector(11 downto 0);
        cd              : out    vl_logic_vector(12 downto 0);
        ctrl            : out    vl_logic_vector(6 downto 0);
        RXen            : out    vl_logic;
        transfer        : out    vl_logic;
        uart_run_flag   : out    vl_logic;
        baud_tick       : out    vl_logic;
        temp_rx_1       : out    vl_logic_vector(11 downto 0);
        rx_fifo_full    : out    vl_logic;
        rx_not_empty    : out    vl_logic;
        rx_write_en     : out    vl_logic;
        rx_read_en      : out    vl_logic;
        data_is_ready   : out    vl_logic;
        rx_ptr_addr_wr_i: out    vl_logic_vector(4 downto 0);
        rx_ptr_addr_rd_o: out    vl_logic_vector(4 downto 0);
        temp_rx         : out    vl_logic_vector(11 downto 0);
        read_data       : out    vl_logic_vector(7 downto 0);
        data_trans      : out    vl_logic_vector(11 downto 0);
        rx_fifo_mid     : out    vl_logic_vector(7 downto 0);
        ctrl_rx_buffer  : out    vl_logic;
        fifo_wr_ctrl    : out    vl_logic;
        data_is_avail   : out    vl_logic;
        RXdone          : out    vl_logic;
        start_bit_rx    : out    vl_logic;
        data_is_received: out    vl_logic;
        parity_bit_rx   : out    vl_logic;
        stop_bit_rx     : out    vl_logic;
        error_rx_detect : out    vl_logic;
        timeout_flag    : out    vl_logic;
        TXdone          : out    vl_logic;
        ctrl_shift_register_rd: out    vl_logic_vector(3 downto 0);
        PREADY          : out    vl_logic;
        PRDATA          : out    vl_logic_vector(31 downto 0)
    );
end test_ver5;
