library verilog;
use verilog.vl_types.all;
entity compare_5bit_vlg_check_tst is
    port(
        A_less_B        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end compare_5bit_vlg_check_tst;
