library verilog;
use verilog.vl_types.all;
entity test_ver5_vlg_vec_tst is
end test_ver5_vlg_vec_tst;
