library verilog;
use verilog.vl_types.all;
entity APB_UART_vlg_vec_tst is
end APB_UART_vlg_vec_tst;
