library verilog;
use verilog.vl_types.all;
entity BAUD_RATE_GENERATOR_vlg_vec_tst is
end BAUD_RATE_GENERATOR_vlg_vec_tst;
