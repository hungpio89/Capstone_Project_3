library verilog;
use verilog.vl_types.all;
entity AHB_APB_UART_vlg_vec_tst is
end AHB_APB_UART_vlg_vec_tst;
