library verilog;
use verilog.vl_types.all;
entity encoder_method_vlg_vec_tst is
end encoder_method_vlg_vec_tst;
