library verilog;
use verilog.vl_types.all;
entity compare_5bit_vlg_vec_tst is
end compare_5bit_vlg_vec_tst;
