library verilog;
use verilog.vl_types.all;
entity ctrl_interface_signal_vlg_vec_tst is
end ctrl_interface_signal_vlg_vec_tst;
