library verilog;
use verilog.vl_types.all;
entity or_1bit_vlg_check_tst is
    port(
        data_out        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end or_1bit_vlg_check_tst;
